class decryptor_configuration extends uvm_object;
	`uvm_object_utils(decryptor_configuration)

	function new(string name = "");
		super.new(name);
	endfunction: new
endclass: decryptor_configuration