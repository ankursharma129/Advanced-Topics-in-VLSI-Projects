// Code your testbench here
// or browse Examples
`include "uvm_macros.svh"
`include "top.sv"
`include "decryptor_bfm.sv"



// `include "scoreboard.svh"
// `include "tester.svh"
// `include "test_bench.svh"
//`include "decryptor_pkg.sv"

