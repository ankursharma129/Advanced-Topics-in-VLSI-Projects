package decryptor_pkg;
import uvm_pkg::*;


	`include "decryptor_sequencer.sv"
	`include "decryptor_monitor.sv"
	`include "decryptor_driver.sv"
	`include "decryptor_agent.sv"
	`include "decryptor_scoreboard.sv"
	`include "decryptor_config.sv"
	`include "decryptor_env.sv"
	`include "decryptor_test.sv"
endpackage : decryptor_pkg