// Code your design here
`include "top_level_4_260.sv"
`include "dat_mem.sv"